module AND_2
(
	input a,b,
	output logic f
);

assign f = a & b;

endmodule: AND_2
