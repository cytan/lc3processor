import lc3b_types::*; /* Import types defined in lc3b_types.sv */

module control
(
    /* Input and output port declarations */
);

enum int unsigned {
    /* List of states */
	 fetch1
} state, next_states;

always_comb
begin : state_actions
    /* Default output assignments */
    /* Actions for each state */
end

always_comb
begin : next_state_logic
    /* Next state information and conditions (if any)
     * for transitioning between states */
end

always_ff @(posedge clk)
begin: next_state_assignment
    /* Assignment of next state on clock edge */
end

endmodule : control
