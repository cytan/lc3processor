module OR_2
(
	input a,b,
	output logic f
);

assign f = a | b;

endmodule: OR_2
